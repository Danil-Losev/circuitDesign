library verilog;
use verilog.vl_types.all;
entity main_vlg_check_tst is
    port(
        F               : in     vl_logic;
        X1              : in     vl_logic;
        X3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end main_vlg_check_tst;
