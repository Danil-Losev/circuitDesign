module main (F, A, B, C); // Определение модуля main с выходом F и входами A, B, C.
    input A, B, C; // Объявление входных сигналов A, B и C.
    output F; // Объявление выходного сигнала F.

    // Присвоение выходу F результата логического выражения:
    // 1. Логическое ИЛИ (OR) между инверсными значениями B и C (~B | ~C).
    // 2. Логическое ИЛИ (OR) между инверсным значением A и B (~A | B).
    // Эти два результата объединяются с помощью логического И (AND).
    assign F = ((~B | ~C) & (~A | B));

endmodule