module main (A, C, G, W); // Определение модуля main с выходом A и входами C, G, W.
    input C, G, W; // Объявление входных сигналов C, G и W.
    output A; // Объявление выходного сигнала A.

    // Присвоение выходу A результата логического выражения, которое состоит из нескольких логических операций:
    // - Логическое И (AND) применяется к результатам нескольких логических ИЛИ (OR):
    //   1. C, G и W
    //   2. C, G и инверсный W
    //   3. C, инверсный G и W
    //   4. Инверсный C, G и W
    //   5. Инверсный C, G и инверсный W
    assign A = ((C|G|W)&(C|G|~W)&(C|~G|W)&(~C|G|W)&(~C|G|~W));

endmodule