library verilog;
use verilog.vl_types.all;
entity main is
    port(
        output_F        : out    vl_logic;
        input_X1        : in     vl_logic;
        input_X3        : in     vl_logic;
        input_X2        : in     vl_logic
    );
end main;
