module main (A, F, C, G, W); // Определение модуля main с выходом A и входами F, C, G, W.
    input F, C, G, W; // Объявление входных сигналов F, C, G и W.
    output A; // Объявление выходного сигнала A.

    // Объявление промежуточных проводов для логических инверсий входных сигналов.
    not(notF, F); // Инвертирование сигнала F, результат сохраняется в notF.
    not(notC, C); // Инвертирование сигнала C, результат сохраняется в notC.
    not(notW, W); // Инвертирование сигнала W, результат сохраняется в notW.
    
    // Логические И для промежуточных сигналов.
    and(and1, notC, W); // AND для инверсного C и W, результат сохраняется в and1.
    and(and2, C, notW); // AND для C и инверсного W, результат сохраняется в and2.
    and(and3, C, W); // AND для C и W, результат сохраняется в and3.

    // Логическое ИЛИ для промежуточных сигналов and1, and2 и and3.
    or(or1, and1, and2, and3); // Результат логического ИЛИ сохраняется в or1.

    // Логическое И для выхода A, использующее G, инверсный F и результат or1.
    and(A, G, notF, or1); // AND для G, notF и or1, результат сохраняется в выходе A.

endmodule