module main (F, A, B, C); // Определение модуля main с выходом F и входами A, B, C.
    input A, B, C; // Объявление входных сигналов A, B и C.
    output F; // Объявление выходного сигнала F.

    // Присвоение выходу F результата логического выражения:
    // 1. Логическое И (AND) между инверсными значениями A и B (~A & ~B).
    // 2. Логическое И (AND) между B и инверсным значением C (B & ~C).
    // Эти два результата объединяются с помощью логического ИЛИ (OR).
    assign F = ((~A & ~B) | (B & ~C));

endmodule