module main (A, C, G, W); // Определение модуля main с входами C, G, W и выходом A.
    input C, G, W; // Объявление входных сигналов C, G и W.
    output A; // Объявление выходного сигнала A.

    wire notC, notG, notW; // Объявление промежуточных проводов для логических инверсий.
    wire temp1, temp2, temp3, temp4, temp5; // Объявление промежуточных проводов для логических операций.

    // Логическое ИЛИ для сигналов C, G и W, результат сохраняется в temp1.
    or(temp1, C, G, W);
    
    // Логическое ИЛИ для сигналов C, G и инверсного W, результат сохраняется в temp2.
    or(temp2, C, G, notW);
    
    // Логическое ИЛИ для сигналов C, инверсного G и W, результат сохраняется в temp3.
    or(temp3, C, notG, W);
    
    // Логическое ИЛИ для инверсного C, G и W, результат сохраняется в temp4.
    or(temp4, notC, G, W);
    
    // Логическое ИЛИ для инверсного C, G и инверсного W, результат сохраняется в temp5.
    or(temp5, notC, G, notW);
    
    // Логическое И AND для всех промежуточных проводов, результат сохраняется в выходе A.
    and(A, temp1, temp2, temp3, temp4, temp5);

endmodule