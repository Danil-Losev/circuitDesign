library verilog;
use verilog.vl_types.all;
entity TaskOneVarSix_vlg_check_tst is
    port(
        output_Y        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TaskOneVarSix_vlg_check_tst;
