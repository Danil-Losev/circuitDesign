module main (F, A, B, C); // Определение модуля main с выходом F и входами A, B, C.
    input A, B, C; // Объявление входных сигналов A, B и C.
    output F; // Объявление выходного сигнала F.

    // Инвертирование входных сигналов A, B и C.
    not(notA, A); // Инвертирование сигнала A, результат сохраняется в notA.
    not(notB, B); // Инвертирование сигнала B, результат сохраняется в notB.
    not(notC, C); // Инвертирование сигнала C, результат сохраняется в notC.

    // Логическое И (AND) для инверсных сигналов A и B.
    and(and1, notA, notB); // AND для notA и notB, результат сохраняется в and1.

    // Логическое И (AND) для сигнала B и инверсного C.
    and(and2, B, notC); // AND для B и notC, результат сохраняется в and2.

    // Логическое ИЛИ (OR) для промежуточных результатов and1 и and2.
    or(F, and1, and2); // OR для and1 и and2, результат сохраняется в выходе F.

endmodule