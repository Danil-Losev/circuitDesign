library verilog;
use verilog.vl_types.all;
entity TaskVar12_vlg_vec_tst is
end TaskVar12_vlg_vec_tst;
