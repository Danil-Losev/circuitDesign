module main (F, A, B, C); // Определение модуля main с выходом F и входами A, B, C.
    input A, B, C; // Объявление входных сигналов A, B и C.
    output F; // Объявление выходного сигнала F.

    // Инвертирование входных сигналов A, B и C.
    not(notA, A); // Инвертирование сигнала A, результат сохраняется в notA.
    not(notB, B); // Инвертирование сигнала B, результат сохраняется в notB.
    not(notC, C); // Инвертирование сигнала C, результат сохраняется в notC.

    // Логическое ИЛИ (OR) для инверсного B и инверсного C.
    or(or1, notB, notC); // OR для notB и notC, результат сохраняется в or1.

    // Логическое ИЛИ (OR) для инверсного A и B.
    or(or2, notA, B); // OR для notA и B, результат сохраняется в or2.

    // Логическое И (AND) для промежуточных результатов or1 и or2.
    and(F, or1, or2); // AND для or1 и or2, результат сохраняется в выходе F.

endmodule