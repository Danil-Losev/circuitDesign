library verilog;
use verilog.vl_types.all;
entity TaskOneVarSix_vlg_vec_tst is
end TaskOneVarSix_vlg_vec_tst;
