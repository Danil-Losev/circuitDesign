library verilog;
use verilog.vl_types.all;
entity TaskVar12_vlg_check_tst is
    port(
        output_F        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TaskVar12_vlg_check_tst;
