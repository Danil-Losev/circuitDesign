library verilog;
use verilog.vl_types.all;
entity TaskVar12 is
    port(
        output_F        : out    vl_logic;
        input_B         : in     vl_logic;
        input_C         : in     vl_logic;
        input_A         : in     vl_logic
    );
end TaskVar12;
