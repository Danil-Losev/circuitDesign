library verilog;
use verilog.vl_types.all;
entity main is
    port(
        F               : out    vl_logic;
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic
    );
end main;
