module main (A, F, C, G, W); // Определение модуля main с выходом A и входами F, C, G, W.
    input F, C, G, W; // Объявление входных сигналов F, C, G и W.
    output A; // Объявление выходного сигнала A.

    // Присвоение выходу A результата логического выражения, которое состоит из:
    // 1. Инверсный сигнал F (~F).
    // 2. Сигнал G.
    // 3. Логическое ИЛИ, состоящее из трех компонентов:
    //    - Инверсный C и W (~C&W).
    //    - C и инверсный W (C&~W).
    //    - C и W (C&W).
    // Все компоненты объединены с помощью логического И (AND).
    assign A = (~F & G & ((~C & W) | (C & ~W) | (C & W))); 

endmodule